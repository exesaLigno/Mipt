module D7seg(input [3:0] dig, output wire [6:0] seg);
    assign seg = (dig==0)? 7'b1000000 :
    (dig==1)? 7'b1111001 :
    (dig==2)? 7'b0100100 :
    (dig==3)? 7'b0110000 :
    (dig==4)? 7'b0011001 :
    (dig==5)? 7'b0010010 :
    (dig==6)? 7'b0000010 :
    (dig==7)? 7'b1111000 :
    (dig==8)? 7'b0000000 :
    (dig==9)? 7'b0010000 :
    (dig=="A")? 7'b1110111 :
    (dig=="b")? 7'b0000011 :
    (dig=="C")? 7'b1000110 :
    (dig=="d")? 7'b0100001 :
    (dig=="E")? 7'b0000110 :
    (dig=="F")? 7'b0001110 :
    7'b1111111 ; // Остальные
endmodule
